magic
tech scmos
timestamp 1731174129
<< nwell >>
rect -7 9 63 94
<< ntransistor >>
rect -6 -24 62 -22
rect -6 -70 62 -68
<< ptransistor >>
rect 22 63 36 65
rect 22 35 36 37
<< ndiffusion >>
rect -6 -12 27 -8
rect 31 -12 62 -8
rect -6 -22 62 -12
rect -6 -38 62 -24
rect -6 -42 27 -38
rect 32 -42 62 -38
rect -6 -58 27 -54
rect 32 -58 62 -54
rect -6 -68 62 -58
rect -6 -84 62 -70
rect -6 -88 27 -84
rect 31 -88 62 -84
<< pdiffusion >>
rect 22 68 26 72
rect 30 68 36 72
rect 22 65 36 68
rect 22 58 36 63
rect 22 54 27 58
rect 32 54 36 58
rect 22 41 27 45
rect 32 41 36 45
rect 22 37 36 41
rect 22 31 36 35
rect 22 27 27 31
rect 31 27 36 31
<< ndcontact >>
rect 27 -12 31 -8
rect 27 -42 32 -38
rect 27 -58 32 -54
rect 27 -88 31 -84
<< pdcontact >>
rect 26 68 30 72
rect 27 54 32 58
rect 27 41 32 45
rect 27 27 31 31
<< psubstratepcontact >>
rect 27 -107 31 -103
rect 37 -107 41 -103
<< nsubstratencontact >>
rect 26 86 30 90
rect 35 86 39 90
<< polysilicon >>
rect -9 63 22 65
rect 36 63 41 65
rect -9 35 22 37
rect 36 35 41 37
rect -7 -24 -6 -22
rect 62 -24 65 -22
rect -9 -70 -6 -68
rect 62 -70 65 -68
<< polycontact >>
rect -14 62 -9 66
rect -13 34 -9 38
rect -11 -25 -7 -21
rect -13 -71 -9 -67
<< metal1 >>
rect -6 86 26 90
rect 30 86 35 90
rect 39 86 62 90
rect 26 72 30 86
rect -23 62 -14 66
rect 27 45 32 54
rect -22 34 -13 38
rect 27 4 31 27
rect 27 -3 88 4
rect 27 -8 31 -3
rect -21 -25 -11 -21
rect 27 -54 32 -42
rect -23 -71 -13 -67
rect 27 -84 31 -83
rect 27 -103 31 -88
rect -23 -107 27 -103
rect 31 -107 37 -103
rect 41 -107 87 -103
rect -23 -109 87 -107
<< labels >>
rlabel metal1 79 1 79 1 1 Vout
rlabel metal1 11 88 11 88 1 Vdd
rlabel metal1 -22 64 -22 64 3 Vbias1
rlabel metal1 -20 36 -20 36 3 Vbias2
rlabel metal1 -19 -23 -19 -23 3 Vbias3
rlabel metal1 -21 -69 -21 -69 3 Vin
<< end >>
