magic
tech scmos
timestamp 1731166859
<< nwell >>
rect -115 -23 158 81
<< ntransistor >>
rect -77 -43 -67 -39
rect -6 -48 14 -44
rect 55 -47 75 -43
rect 130 -46 150 -42
rect -6 -92 14 -88
rect 56 -91 76 -87
rect 131 -93 151 -89
<< ptransistor >>
rect 101 42 149 46
rect -82 -1 -34 3
rect -19 -1 29 3
rect 45 -1 85 9
rect 101 -1 149 3
<< ndiffusion >>
rect -77 -35 -74 -31
rect -70 -35 -67 -31
rect -77 -39 -67 -35
rect -6 -41 -1 -37
rect 3 -41 14 -37
rect -77 -45 -67 -43
rect -6 -44 14 -41
rect 55 -40 62 -36
rect 66 -40 75 -36
rect 55 -43 75 -40
rect 130 -39 136 -35
rect 140 -39 150 -35
rect 130 -42 150 -39
rect -77 -49 -76 -45
rect -72 -49 -67 -45
rect -77 -50 -67 -49
rect -6 -51 14 -48
rect -6 -55 -1 -51
rect 3 -55 14 -51
rect 55 -50 75 -47
rect 55 -54 62 -50
rect 66 -54 75 -50
rect 130 -49 150 -46
rect 130 -53 136 -49
rect 140 -53 150 -49
rect -6 -86 -1 -82
rect 3 -86 14 -82
rect -6 -88 14 -86
rect 56 -85 62 -81
rect 66 -85 76 -81
rect 56 -87 76 -85
rect 131 -87 136 -83
rect 140 -87 151 -83
rect 131 -89 151 -87
rect -6 -94 14 -92
rect -6 -98 -4 -94
rect 0 -98 14 -94
rect 56 -93 76 -91
rect 56 -97 57 -93
rect 61 -97 76 -93
rect 131 -95 151 -93
rect 131 -99 133 -95
rect 137 -99 151 -95
<< pdiffusion >>
rect 101 56 149 57
rect 101 52 103 56
rect 107 52 149 56
rect 101 46 149 52
rect 101 38 149 42
rect 101 34 121 38
rect 125 34 149 38
rect 101 31 149 34
rect -82 10 -77 14
rect -73 10 -34 14
rect -82 3 -34 10
rect -19 13 29 14
rect -19 9 -13 13
rect -9 9 29 13
rect 45 11 48 15
rect 52 11 85 15
rect 45 9 85 11
rect 101 12 149 14
rect -19 3 29 9
rect 101 8 121 12
rect 125 8 149 12
rect 101 3 149 8
rect -82 -8 -34 -1
rect -82 -12 -74 -8
rect -70 -12 -34 -8
rect -19 -7 29 -1
rect -19 -11 -1 -7
rect 3 -11 29 -7
rect -19 -12 29 -11
rect 45 -7 85 -1
rect 45 -11 62 -7
rect 66 -11 85 -7
rect 45 -12 85 -11
rect 101 -7 149 -1
rect 101 -11 136 -7
rect 140 -11 149 -7
rect 101 -12 149 -11
<< ndcontact >>
rect -74 -35 -70 -31
rect -1 -41 3 -37
rect 62 -40 66 -36
rect 136 -39 140 -35
rect -76 -49 -72 -45
rect -1 -55 3 -51
rect 62 -54 66 -50
rect 136 -53 140 -49
rect -1 -86 3 -82
rect 62 -85 66 -81
rect 136 -87 140 -83
rect -4 -98 0 -94
rect 57 -97 61 -93
rect 133 -99 137 -95
<< pdcontact >>
rect 103 52 107 56
rect 121 34 125 38
rect -77 10 -73 14
rect -13 9 -9 13
rect 48 11 52 15
rect 121 8 125 12
rect -74 -12 -70 -8
rect -1 -11 3 -7
rect 62 -11 66 -7
rect 136 -11 140 -7
<< psubstratepcontact >>
rect -76 -108 -72 -104
rect -67 -108 -63 -104
rect -4 -108 0 -104
rect 4 -108 8 -104
rect 57 -108 61 -104
rect 66 -108 70 -104
rect 133 -108 137 -104
rect 142 -108 146 -104
<< nsubstratencontact >>
rect -77 72 -73 76
rect -66 72 -62 76
rect -13 71 -9 75
rect -4 71 0 75
rect 48 71 52 75
rect 56 71 60 75
rect 103 71 107 75
rect 111 71 115 75
<< polysilicon >>
rect 98 42 101 46
rect 149 42 151 46
rect -85 -1 -82 3
rect -34 -1 -19 3
rect 29 -1 33 3
rect 36 -1 45 9
rect 85 -1 90 9
rect 94 -1 101 3
rect 149 -1 151 3
rect -85 -43 -77 -39
rect -67 -43 -64 -39
rect 43 -44 55 -43
rect -7 -48 -6 -44
rect 14 -47 55 -44
rect 75 -47 76 -43
rect 128 -46 130 -42
rect 150 -46 155 -42
rect 14 -48 43 -47
rect -12 -92 -6 -88
rect 14 -92 16 -88
rect 53 -91 56 -87
rect 76 -91 78 -87
rect 129 -93 131 -89
rect 151 -93 155 -89
<< polycontact >>
rect 151 42 155 46
rect -89 -1 -85 3
rect 90 -1 94 3
rect 151 -1 155 3
rect -64 -43 -60 -39
rect -11 -48 -7 -44
rect 76 -47 80 -43
rect 124 -46 128 -42
rect 16 -92 20 -88
rect 49 -91 53 -87
rect 78 -91 82 -87
rect 125 -93 129 -89
<< metal1 >>
rect -87 76 148 79
rect -87 72 -77 76
rect -73 72 -66 76
rect -62 75 148 76
rect -62 72 -13 75
rect -87 71 -13 72
rect -9 71 -4 75
rect 0 71 48 75
rect 52 71 56 75
rect 60 71 103 75
rect 107 71 111 75
rect 115 71 148 75
rect -87 70 148 71
rect -77 14 -73 70
rect -13 13 -9 70
rect 48 15 52 70
rect 103 56 107 70
rect 155 42 165 46
rect 121 38 125 40
rect 121 12 125 34
rect 121 6 125 8
rect 159 11 163 42
rect 159 7 177 11
rect -100 -1 -89 3
rect 155 -1 159 3
rect -74 -27 -70 -12
rect -74 -30 -51 -27
rect -74 -31 -70 -30
rect -74 -36 -70 -35
rect -55 -39 -51 -30
rect -1 -31 3 -11
rect 62 -18 66 -11
rect 90 -18 94 -1
rect 173 -5 177 7
rect 62 -22 94 -18
rect 136 -7 140 -6
rect 136 -18 140 -11
rect 159 -9 177 -5
rect 159 -18 163 -9
rect 136 -22 163 -18
rect -1 -35 28 -31
rect -1 -37 3 -35
rect -60 -43 -20 -39
rect -25 -44 -20 -43
rect 24 -44 28 -35
rect 62 -36 66 -22
rect 136 -35 140 -22
rect 136 -40 140 -39
rect 62 -41 66 -40
rect 118 -43 124 -42
rect -25 -48 -11 -44
rect 80 -46 124 -43
rect 80 -47 122 -46
rect -76 -103 -72 -49
rect -1 -82 3 -55
rect 24 -88 28 -48
rect 62 -81 66 -54
rect 136 -83 140 -53
rect 40 -88 49 -87
rect 20 -91 49 -88
rect 82 -89 104 -87
rect 82 -91 125 -89
rect 20 -92 44 -91
rect 100 -93 125 -91
rect -4 -103 0 -98
rect 57 -103 61 -97
rect 133 -103 137 -99
rect -110 -104 185 -103
rect -110 -108 -76 -104
rect -72 -108 -67 -104
rect -63 -108 -4 -104
rect 0 -108 4 -104
rect 8 -108 57 -104
rect 61 -108 66 -104
rect 70 -108 133 -104
rect 137 -108 142 -104
rect 146 -108 185 -104
rect -110 -112 185 -108
<< labels >>
rlabel metal1 28 -108 28 -108 1 gnd!
rlabel metal1 -100 -1 -100 3 1 vin
rlabel metal1 -56 74 -56 74 1 vdd
rlabel metal1 165 42 165 46 1 vbias1
rlabel metal1 159 -1 159 3 1 vbias2
<< end >>
